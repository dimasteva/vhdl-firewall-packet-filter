LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE std.textio.ALL;

-- WHEN RUNNING THE TESTBENCH IT WILL END WITH THE MESSAGE END
-- AFTER THAT MESSAGE IT WILL SAY 'REPORT FAILED' AND 'SIMULATION FAILED' BUT PAY NO MIND TO THAT

-- EVERY TIME THE OUT_WRITE_ENABLE SIGNAL IS SET THE TESTBENCH WILL PRINT THE OUTPUT
-- TO THE CONSOLE INSTEAD OF WRITING IT INTO THE MEMORY

-- IT _MAY_ HAVE BUGS :)


ENTITY project_io_tb IS
GENERIC (
    IN_RAM_SIZE : NATURAL := 1500;
    OUT_RAM_SIZE : NATURAL := 2;
    BUFFER_NUM : NATURAL := 1
);
END ENTITY project_io_tb;

ARCHITECTURE behavioural OF project_io_tb IS
    COMPONENT project_io IS
        PORT (
            clk : IN STD_LOGIC;
            rst : IN STD_LOGIC;
            enable : IN STD_LOGIC;
            done : OUT STD_LOGIC;
            in_read_enable : OUT STD_LOGIC;
            in_index : OUT INTEGER;
            in_data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
            out_write_enable : OUT STD_LOGIC;
            out_index : OUT INTEGER;
            out_data : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
            in_buff_size : OUT INTEGER;
            out_buff_size : OUT INTEGER
        );
    END COMPONENT;
    
    TYPE memory_array IS ARRAY(natural RANGE <>) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE memory_bank IS ARRAY(natural RANGE <>) OF memory_array(0 to IN_RAM_SIZE-1);
    -- RAM
    SIGNAL in_ram : memory_array (0 TO IN_RAM_SIZE-1);
    SIGNAL out_ram : memory_array (0 TO OUT_RAM_SIZE-1);

    -- SIGNALS IN PROJECT_IO
    SIGNAL clk : STD_LOGIC;
    SIGNAL rst : STD_LOGIC := '0';
    SIGNAL enable : STD_LOGIC := '0';
    SIGNAL in_data : STD_LOGIC_VECTOR(7 DOWNTO 0);

    -- SIGNALS OUT PROJECT_IO
    SIGNAL done : STD_LOGIC;
    SIGNAL in_read_enable : STD_LOGIC;
    SIGNAL in_index : INTEGER;
    SIGNAL out_write_enable : STD_LOGIC;
    SIGNAL out_index : INTEGER;
    SIGNAL out_data : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL in_buff_size : INTEGER;
    SIGNAL out_buff_size : INTEGER;

    -- INTERNAL SIGNALS
    SIGNAL curr_buffer : INTEGER := 0;


    -- THIS IS WHERE YOU PUT YOUR BUFFERS
    -- AFTER EVERY GIVEN ONE TACT SIGNAL 'DONE' THE NEXT BUFFER IS LOADED
    SIGNAL buffer_array : memory_bank (0 to BUFFER_NUM-1) := (
    0 => (
        0 => X"00", 1 => X"00",
        2 => X"00", 3 => X"01",
        4 => X"00", 5 => X"02",
        6 => X"00", 7 => X"03",
        8 => X"00", 9 => X"04",
        10 => X"00", 11 => X"05",
        12 => X"00", 13 => X"06",
        14 => X"00", 15 => X"07",
        16 => X"00", 17 => X"08",
        18 => X"00", 19 => X"09",
        20 => X"00", 21 => X"0A",
        22 => X"00", 23 => X"0B",
        24 => X"00", 25 => X"0C",
        26 => X"00", 27 => X"0D",
        28 => X"00", 29 => X"0E",
        30 => X"00", 31 => X"0F",
        32 => X"00", 33 => X"10",
        34 => X"00", 35 => X"11",
        36 => X"00", 37 => X"12",
        38 => X"00", 39 => X"13",
        40 => X"00", 41 => X"14",
        42 => X"00", 43 => X"15",
        44 => X"00", 45 => X"16",
        46 => X"00", 47 => X"17",
        48 => X"00", 49 => X"18",
        50 => X"00", 51 => X"19",
        52 => X"00", 53 => X"1A",
        54 => X"00", 55 => X"1B",
        56 => X"00", 57 => X"1C",
        58 => X"00", 59 => X"1D",
        60 => X"00", 61 => X"1E",
        62 => X"00", 63 => X"1F",
        64 => X"00", 65 => X"20",
        66 => X"00", 67 => X"21",
        68 => X"00", 69 => X"22",
        70 => X"00", 71 => X"23",
        72 => X"00", 73 => X"24",
        74 => X"00", 75 => X"25",
        76 => X"00", 77 => X"26",
        78 => X"00", 79 => X"27",
        80 => X"00", 81 => X"28",
        82 => X"00", 83 => X"29",
        84 => X"00", 85 => X"2A",
        86 => X"00", 87 => X"2B",
        88 => X"00", 89 => X"2C",
        90 => X"00", 91 => X"2D",
        92 => X"00", 93 => X"2E",
        94 => X"00", 95 => X"2F",
        96 => X"00", 97 => X"30",
        98 => X"00", 99 => X"31",
        100 => X"00", 101 => X"32",
        102 => X"00", 103 => X"33",
        104 => X"00", 105 => X"34",
        106 => X"00", 107 => X"35",
        108 => X"00", 109 => X"36",
        110 => X"00", 111 => X"37",
        112 => X"00", 113 => X"38",
        114 => X"00", 115 => X"39",
        116 => X"00", 117 => X"3A",
        118 => X"00", 119 => X"3B",
        120 => X"00", 121 => X"3C",
        122 => X"00", 123 => X"3D",
        124 => X"00", 125 => X"3E",
        126 => X"00", 127 => X"3F",
        128 => X"00", 129 => X"40",
        130 => X"00", 131 => X"41",
        132 => X"00", 133 => X"42",
        134 => X"00", 135 => X"43",
        136 => X"00", 137 => X"44",
        138 => X"00", 139 => X"45",
        140 => X"00", 141 => X"46",
        142 => X"00", 143 => X"47",
        144 => X"00", 145 => X"48",
        146 => X"00", 147 => X"49",
        148 => X"00", 149 => X"4A",
        150 => X"00", 151 => X"4B",
        152 => X"00", 153 => X"4C",
        154 => X"00", 155 => X"4D",
        156 => X"00", 157 => X"4E",
        158 => X"00", 159 => X"4F",
        160 => X"00", 161 => X"50",
        162 => X"00", 163 => X"51",
        164 => X"00", 165 => X"52",
        166 => X"00", 167 => X"53",
        168 => X"00", 169 => X"54",
        170 => X"00", 171 => X"55",
        172 => X"00", 173 => X"56",
        174 => X"00", 175 => X"57",
        176 => X"00", 177 => X"58",
        178 => X"00", 179 => X"59",
        180 => X"00", 181 => X"5A",
        182 => X"00", 183 => X"5B",
        184 => X"00", 185 => X"5C",
        186 => X"00", 187 => X"5D",
        188 => X"00", 189 => X"5E",
        190 => X"00", 191 => X"5F",
        192 => X"00", 193 => X"60",
        194 => X"00", 195 => X"61",
        196 => X"00", 197 => X"62",
        198 => X"00", 199 => X"63",
        200 => X"00", 201 => X"64",
        202 => X"00", 203 => X"65",
        204 => X"00", 205 => X"66",
        206 => X"00", 207 => X"67",
        208 => X"00", 209 => X"68",
        210 => X"00", 211 => X"69",
        212 => X"00", 213 => X"6A",
        214 => X"00", 215 => X"6B",
        216 => X"00", 217 => X"6C",
        218 => X"00", 219 => X"6D",
        220 => X"00", 221 => X"6E",
        222 => X"00", 223 => X"6F",
        224 => X"00", 225 => X"70",
        226 => X"00", 227 => X"71",
        228 => X"00", 229 => X"72",
        230 => X"00", 231 => X"73",
        232 => X"00", 233 => X"74",
        234 => X"00", 235 => X"75",
        236 => X"00", 237 => X"76",
        238 => X"00", 239 => X"77",
        240 => X"00", 241 => X"78",
        242 => X"00", 243 => X"79",
        244 => X"00", 245 => X"7A",
        246 => X"00", 247 => X"7B",
        248 => X"00", 249 => X"7C",
        250 => X"00", 251 => X"7D",
        252 => X"00", 253 => X"7E",
        254 => X"00", 255 => X"7F",
        256 => X"00", 257 => X"80",
        258 => X"00", 259 => X"81",
        260 => X"00", 261 => X"82",
        262 => X"00", 263 => X"83",
        264 => X"00", 265 => X"84",
        266 => X"00", 267 => X"85",
        268 => X"00", 269 => X"86",
        270 => X"00", 271 => X"87",
        272 => X"00", 273 => X"88",
        274 => X"00", 275 => X"89",
        276 => X"00", 277 => X"8A",
        278 => X"00", 279 => X"8B",
        280 => X"00", 281 => X"8C",
        282 => X"00", 283 => X"8D",
        284 => X"00", 285 => X"8E",
        286 => X"00", 287 => X"8F",
        288 => X"00", 289 => X"90",
        290 => X"00", 291 => X"91",
        292 => X"00", 293 => X"92",
        294 => X"00", 295 => X"93",
        296 => X"00", 297 => X"94",
        298 => X"00", 299 => X"95",
        300 => X"00", 301 => X"96",
        302 => X"00", 303 => X"97",
        304 => X"00", 305 => X"98",
        306 => X"00", 307 => X"99",
        308 => X"00", 309 => X"9A",
        310 => X"00", 311 => X"9B",
        312 => X"00", 313 => X"9C",
        314 => X"00", 315 => X"9D",
        316 => X"00", 317 => X"9E",
        318 => X"00", 319 => X"9F",
        320 => X"00", 321 => X"A0",
        322 => X"00", 323 => X"A1",
        324 => X"00", 325 => X"A2",
        326 => X"00", 327 => X"A3",
        328 => X"00", 329 => X"A4",
        330 => X"00", 331 => X"A5",
        332 => X"00", 333 => X"A6",
        334 => X"00", 335 => X"A7",
        336 => X"00", 337 => X"A8",
        338 => X"00", 339 => X"A9",
        340 => X"00", 341 => X"AA",
        342 => X"00", 343 => X"AB",
        344 => X"00", 345 => X"AC",
        346 => X"00", 347 => X"AD",
        348 => X"00", 349 => X"AE",
        350 => X"00", 351 => X"AF",
        352 => X"00", 353 => X"B0",
        354 => X"00", 355 => X"B1",
        356 => X"00", 357 => X"B2",
        358 => X"00", 359 => X"B3",
        360 => X"00", 361 => X"B4",
        362 => X"00", 363 => X"B5",
        364 => X"00", 365 => X"B6",
        366 => X"00", 367 => X"B7",
        368 => X"00", 369 => X"B8",
        370 => X"00", 371 => X"B9",
        372 => X"00", 373 => X"BA",
        374 => X"00", 375 => X"BB",
        376 => X"00", 377 => X"BC",
        378 => X"00", 379 => X"BD",
        380 => X"00", 381 => X"BE",
        382 => X"00", 383 => X"BF",
        384 => X"00", 385 => X"C0",
        386 => X"00", 387 => X"C1",
        388 => X"00", 389 => X"C2",
        390 => X"00", 391 => X"C3",
        392 => X"00", 393 => X"C4",
        394 => X"00", 395 => X"C5",
        396 => X"00", 397 => X"C6",
        398 => X"00", 399 => X"C7",
        400 => X"00", 401 => X"C8",
        402 => X"00", 403 => X"C9",
        404 => X"00", 405 => X"CA",
        406 => X"00", 407 => X"CB",
        408 => X"00", 409 => X"CC",
        410 => X"00", 411 => X"CD",
        412 => X"00", 413 => X"CE",
        414 => X"00", 415 => X"CF",
        416 => X"00", 417 => X"D0",
        418 => X"00", 419 => X"D1",
        420 => X"00", 421 => X"D2",
        422 => X"00", 423 => X"D3",
        424 => X"00", 425 => X"D4",
        426 => X"00", 427 => X"D5",
        428 => X"00", 429 => X"D6",
        430 => X"00", 431 => X"D7",
        432 => X"00", 433 => X"D8",
        434 => X"00", 435 => X"D9",
        436 => X"00", 437 => X"DA",
        438 => X"00", 439 => X"DB",
        440 => X"00", 441 => X"DC",
        442 => X"00", 443 => X"DD",
        444 => X"00", 445 => X"DE",
        446 => X"00", 447 => X"DF",
        448 => X"00", 449 => X"E0",
        450 => X"00", 451 => X"E1",
        452 => X"00", 453 => X"E2",
        454 => X"00", 455 => X"E3",
        456 => X"00", 457 => X"E4",
        458 => X"00", 459 => X"E5",
        460 => X"00", 461 => X"E6",
        462 => X"00", 463 => X"E7",
        464 => X"00", 465 => X"E8",
        466 => X"00", 467 => X"E9",
        468 => X"00", 469 => X"EA",
        470 => X"00", 471 => X"EB",
        472 => X"00", 473 => X"EC",
        474 => X"00", 475 => X"ED",
        476 => X"00", 477 => X"EE",
        478 => X"00", 479 => X"EF",
        480 => X"00", 481 => X"F0",
        482 => X"00", 483 => X"F1",
        484 => X"00", 485 => X"F2",
        486 => X"00", 487 => X"F3",
        488 => X"00", 489 => X"F4",
        490 => X"00", 491 => X"F5",
        492 => X"00", 493 => X"F6",
        494 => X"00", 495 => X"F7",
        496 => X"00", 497 => X"F8",
        498 => X"00", 499 => X"F9",
        500 => X"00", 501 => X"FA",
        502 => X"00", 503 => X"FB",
        504 => X"00", 505 => X"FC",
        506 => X"00", 507 => X"FD",
        508 => X"00", 509 => X"FE",
        510 => X"00", 511 => X"FF",
        512 => X"01", 513 => X"00",
        514 => X"01", 515 => X"01",
        516 => X"01", 517 => X"02",
        518 => X"01", 519 => X"03",
        520 => X"01", 521 => X"04",
        522 => X"01", 523 => X"05",
        524 => X"01", 525 => X"06",
        526 => X"01", 527 => X"07",
        528 => X"01", 529 => X"08",
        530 => X"01", 531 => X"09",
        532 => X"01", 533 => X"0A",
        534 => X"01", 535 => X"0B",
        536 => X"01", 537 => X"0C",
        538 => X"01", 539 => X"0D",
        540 => X"01", 541 => X"0E",
        542 => X"01", 543 => X"0F",
        544 => X"01", 545 => X"10",
        546 => X"01", 547 => X"11",
        548 => X"01", 549 => X"12",
        550 => X"01", 551 => X"13",
        552 => X"01", 553 => X"14",
        554 => X"01", 555 => X"15",
        556 => X"01", 557 => X"16",
        558 => X"01", 559 => X"17",
        560 => X"01", 561 => X"18",
        562 => X"01", 563 => X"19",
        564 => X"01", 565 => X"1A",
        566 => X"01", 567 => X"1B",
        568 => X"01", 569 => X"1C",
        570 => X"01", 571 => X"1D",
        572 => X"01", 573 => X"1E",
        574 => X"01", 575 => X"1F",
        576 => X"01", 577 => X"20",
        578 => X"01", 579 => X"21",
        580 => X"01", 581 => X"22",
        582 => X"01", 583 => X"23",
        584 => X"01", 585 => X"24",
        586 => X"01", 587 => X"25",
        588 => X"01", 589 => X"26",
        590 => X"01", 591 => X"27",
        592 => X"01", 593 => X"28",
        594 => X"01", 595 => X"29",
        596 => X"01", 597 => X"2A",
        598 => X"01", 599 => X"2B",
        600 => X"01", 601 => X"2C",
        602 => X"01", 603 => X"2D",
        604 => X"01", 605 => X"2E",
        606 => X"01", 607 => X"2F",
        608 => X"01", 609 => X"30",
        610 => X"01", 611 => X"31",
        612 => X"01", 613 => X"32",
        614 => X"01", 615 => X"33",
        616 => X"01", 617 => X"34",
        618 => X"01", 619 => X"35",
        620 => X"01", 621 => X"36",
        622 => X"01", 623 => X"37",
        624 => X"01", 625 => X"38",
        626 => X"01", 627 => X"39",
        628 => X"01", 629 => X"3A",
        630 => X"01", 631 => X"3B",
        632 => X"01", 633 => X"3C",
        634 => X"01", 635 => X"3D",
        636 => X"01", 637 => X"3E",
        638 => X"01", 639 => X"3F",
        640 => X"01", 641 => X"40",
        642 => X"01", 643 => X"41",
        644 => X"01", 645 => X"42",
        646 => X"01", 647 => X"43",
        648 => X"01", 649 => X"44",
        650 => X"01", 651 => X"45",
        652 => X"01", 653 => X"46",
        654 => X"01", 655 => X"47",
        656 => X"01", 657 => X"48",
        658 => X"01", 659 => X"49",
        660 => X"01", 661 => X"4A",
        662 => X"01", 663 => X"4B",
        664 => X"01", 665 => X"4C",
        666 => X"01", 667 => X"4D",
        668 => X"01", 669 => X"4E",
        670 => X"01", 671 => X"4F",
        672 => X"01", 673 => X"50",
        674 => X"01", 675 => X"51",
        676 => X"01", 677 => X"52",
        678 => X"01", 679 => X"53",
        680 => X"01", 681 => X"54",
        682 => X"01", 683 => X"55",
        684 => X"01", 685 => X"56",
        686 => X"01", 687 => X"57",
        688 => X"01", 689 => X"58",
        690 => X"01", 691 => X"59",
        692 => X"01", 693 => X"5A",
        694 => X"01", 695 => X"5B",
        696 => X"01", 697 => X"5C",
        698 => X"01", 699 => X"5D",
        700 => X"01", 701 => X"5E",
        702 => X"01", 703 => X"5F",
        704 => X"01", 705 => X"60",
        706 => X"01", 707 => X"61",
        708 => X"01", 709 => X"62",
        710 => X"01", 711 => X"63",
        712 => X"01", 713 => X"64",
        714 => X"01", 715 => X"65",
        716 => X"01", 717 => X"66",
        718 => X"01", 719 => X"67",
        720 => X"01", 721 => X"68",
        722 => X"01", 723 => X"69",
        724 => X"01", 725 => X"6A",
        726 => X"01", 727 => X"6B",
        728 => X"01", 729 => X"6C",
        730 => X"01", 731 => X"6D",
        732 => X"01", 733 => X"6E",
        734 => X"01", 735 => X"6F",
        736 => X"01", 737 => X"70",
        738 => X"01", 739 => X"71",
        740 => X"01", 741 => X"72",
        742 => X"01", 743 => X"73",
        744 => X"01", 745 => X"74",
        746 => X"01", 747 => X"75",
        748 => X"01", 749 => X"76",
        750 => X"01", 751 => X"77",
        752 => X"01", 753 => X"78",
        754 => X"01", 755 => X"79",
        756 => X"01", 757 => X"7A",
        758 => X"01", 759 => X"7B",
        760 => X"01", 761 => X"7C",
        762 => X"01", 763 => X"7D",
        764 => X"01", 765 => X"7E",
        766 => X"01", 767 => X"7F",
        768 => X"01", 769 => X"80",
        770 => X"01", 771 => X"81",
        772 => X"01", 773 => X"82",
        774 => X"01", 775 => X"83",
        776 => X"01", 777 => X"84",
        778 => X"01", 779 => X"85",
        780 => X"01", 781 => X"86",
        782 => X"01", 783 => X"87",
        784 => X"01", 785 => X"88",
        786 => X"01", 787 => X"89",
        788 => X"01", 789 => X"8A",
        790 => X"01", 791 => X"8B",
        792 => X"01", 793 => X"8C",
        794 => X"01", 795 => X"8D",
        796 => X"01", 797 => X"8E",
        798 => X"01", 799 => X"8F",
        800 => X"01", 801 => X"90",
        802 => X"01", 803 => X"91",
        804 => X"01", 805 => X"92",
        806 => X"01", 807 => X"93",
        808 => X"01", 809 => X"94",
        810 => X"01", 811 => X"95",
        812 => X"01", 813 => X"96",
        814 => X"01", 815 => X"97",
        816 => X"01", 817 => X"98",
        818 => X"01", 819 => X"99",
        820 => X"01", 821 => X"9A",
        822 => X"01", 823 => X"9B",
        824 => X"01", 825 => X"9C",
        826 => X"01", 827 => X"9D",
        828 => X"01", 829 => X"9E",
        830 => X"01", 831 => X"9F",
        832 => X"01", 833 => X"A0",
        834 => X"01", 835 => X"A1",
        836 => X"01", 837 => X"A2",
        838 => X"01", 839 => X"A3",
        840 => X"01", 841 => X"A4",
        842 => X"01", 843 => X"A5",
        844 => X"01", 845 => X"A6",
        846 => X"01", 847 => X"A7",
        848 => X"01", 849 => X"A8",
        850 => X"01", 851 => X"A9",
        852 => X"01", 853 => X"AA",
        854 => X"01", 855 => X"AB",
        856 => X"01", 857 => X"AC",
        858 => X"01", 859 => X"AD",
        860 => X"01", 861 => X"AE",
        862 => X"01", 863 => X"AF",
        864 => X"01", 865 => X"B0",
        866 => X"01", 867 => X"B1",
        868 => X"01", 869 => X"B2",
        870 => X"01", 871 => X"B3",
        872 => X"01", 873 => X"B4",
        874 => X"01", 875 => X"B5",
        876 => X"01", 877 => X"B6",
        878 => X"01", 879 => X"B7",
        880 => X"01", 881 => X"B8",
        882 => X"01", 883 => X"B9",
        884 => X"01", 885 => X"BA",
        886 => X"01", 887 => X"BB",
        888 => X"01", 889 => X"BC",
        890 => X"01", 891 => X"BD",
        892 => X"01", 893 => X"BE",
        894 => X"01", 895 => X"BF",
        896 => X"01", 897 => X"C0",
        898 => X"01", 899 => X"C1",
        900 => X"01", 901 => X"C2",
        902 => X"01", 903 => X"C3",
        904 => X"01", 905 => X"C4",
        906 => X"01", 907 => X"C5",
        908 => X"01", 909 => X"C6",
        910 => X"01", 911 => X"C7",
        912 => X"01", 913 => X"C8",
        914 => X"01", 915 => X"C9",
        916 => X"01", 917 => X"CA",
        918 => X"01", 919 => X"CB",
        920 => X"01", 921 => X"CC",
        922 => X"01", 923 => X"CD",
        924 => X"01", 925 => X"CE",
        926 => X"01", 927 => X"CF",
        928 => X"01", 929 => X"D0",
        930 => X"01", 931 => X"D1",
        932 => X"01", 933 => X"D2",
        934 => X"01", 935 => X"D3",
        936 => X"01", 937 => X"D4",
        938 => X"01", 939 => X"D5",
        940 => X"01", 941 => X"D6",
        942 => X"01", 943 => X"D7",
        944 => X"01", 945 => X"D8",
        946 => X"01", 947 => X"D9",
        948 => X"01", 949 => X"DA",
        950 => X"01", 951 => X"DB",
        952 => X"01", 953 => X"DC",
        954 => X"01", 955 => X"DD",
        956 => X"01", 957 => X"DE",
        958 => X"01", 959 => X"DF",
        960 => X"01", 961 => X"E0",
        962 => X"01", 963 => X"E1",
        964 => X"01", 965 => X"E2",
        966 => X"01", 967 => X"E3",
        968 => X"01", 969 => X"E4",
        970 => X"01", 971 => X"E5",
        972 => X"01", 973 => X"E6",
        974 => X"01", 975 => X"E7",
        976 => X"01", 977 => X"E8",
        978 => X"01", 979 => X"E9",
        980 => X"01", 981 => X"EA",
        982 => X"01", 983 => X"EB",
        984 => X"01", 985 => X"EC",
        986 => X"01", 987 => X"ED",
        988 => X"01", 989 => X"EE",
        990 => X"01", 991 => X"EF",
        992 => X"01", 993 => X"F0",
        994 => X"01", 995 => X"F1",
        996 => X"01", 997 => X"F2",
        998 => X"01", 999 => X"F3",
        1000 => X"01", 1001 => X"F4",
        1002 => X"01", 1003 => X"F5",
        1004 => X"01", 1005 => X"F6",
        1006 => X"01", 1007 => X"F7",
        1008 => X"01", 1009 => X"F8",
        1010 => X"01", 1011 => X"F9",
        1012 => X"01", 1013 => X"FA",
        1014 => X"01", 1015 => X"FB",
        1016 => X"01", 1017 => X"FC",
        1018 => X"01", 1019 => X"FD",
        1020 => X"01", 1021 => X"FE",
        1022 => X"01", 1023 => X"FF",
        1024 => X"02", 1025 => X"00",
        1026 => X"02", 1027 => X"01",
        1028 => X"02", 1029 => X"02",
        1030 => X"02", 1031 => X"03",
        1032 => X"02", 1033 => X"04",
        1034 => X"02", 1035 => X"05",
        1036 => X"02", 1037 => X"06",
        1038 => X"02", 1039 => X"07",
        1040 => X"02", 1041 => X"08",
        1042 => X"02", 1043 => X"09",
        1044 => X"02", 1045 => X"0A",
        1046 => X"02", 1047 => X"0B",
        1048 => X"02", 1049 => X"0C",
        1050 => X"02", 1051 => X"0D",
        1052 => X"02", 1053 => X"0E",
        1054 => X"02", 1055 => X"0F",
        1056 => X"02", 1057 => X"10",
        1058 => X"02", 1059 => X"11",
        1060 => X"02", 1061 => X"12",
        1062 => X"02", 1063 => X"13",
        1064 => X"02", 1065 => X"14",
        1066 => X"02", 1067 => X"15",
        1068 => X"02", 1069 => X"16",
        1070 => X"02", 1071 => X"17",
        1072 => X"02", 1073 => X"18",
        1074 => X"02", 1075 => X"19",
        1076 => X"02", 1077 => X"1A",
        1078 => X"02", 1079 => X"1B",
        1080 => X"02", 1081 => X"1C",
        1082 => X"02", 1083 => X"1D",
        1084 => X"02", 1085 => X"1E",
        1086 => X"02", 1087 => X"1F",
        1088 => X"02", 1089 => X"20",
        1090 => X"02", 1091 => X"21",
        1092 => X"02", 1093 => X"22",
        1094 => X"02", 1095 => X"23",
        1096 => X"02", 1097 => X"24",
        1098 => X"02", 1099 => X"25",
        1100 => X"02", 1101 => X"26",
        1102 => X"02", 1103 => X"27",
        1104 => X"02", 1105 => X"28",
        1106 => X"02", 1107 => X"29",
        1108 => X"02", 1109 => X"2A",
        1110 => X"02", 1111 => X"2B",
        1112 => X"02", 1113 => X"2C",
        1114 => X"02", 1115 => X"2D",
        1116 => X"02", 1117 => X"2E",
        1118 => X"02", 1119 => X"2F",
        1120 => X"02", 1121 => X"30",
        1122 => X"02", 1123 => X"31",
        1124 => X"02", 1125 => X"32",
        1126 => X"02", 1127 => X"33",
        1128 => X"02", 1129 => X"34",
        1130 => X"02", 1131 => X"35",
        1132 => X"02", 1133 => X"36",
        1134 => X"02", 1135 => X"37",
        1136 => X"02", 1137 => X"38",
        1138 => X"02", 1139 => X"39",
        1140 => X"02", 1141 => X"3A",
        1142 => X"02", 1143 => X"3B",
        1144 => X"02", 1145 => X"3C",
        1146 => X"02", 1147 => X"3D",
        1148 => X"02", 1149 => X"3E",
        1150 => X"02", 1151 => X"3F",
        1152 => X"02", 1153 => X"40",
        1154 => X"02", 1155 => X"41",
        1156 => X"02", 1157 => X"42",
        1158 => X"02", 1159 => X"43",
        1160 => X"02", 1161 => X"44",
        1162 => X"02", 1163 => X"45",
        1164 => X"02", 1165 => X"46",
        1166 => X"02", 1167 => X"47",
        1168 => X"02", 1169 => X"48",
        1170 => X"02", 1171 => X"49",
        1172 => X"02", 1173 => X"4A",
        1174 => X"02", 1175 => X"4B",
        1176 => X"02", 1177 => X"4C",
        1178 => X"02", 1179 => X"4D",
        1180 => X"02", 1181 => X"4E",
        1182 => X"02", 1183 => X"4F",
        1184 => X"02", 1185 => X"50",
        1186 => X"02", 1187 => X"51",
        1188 => X"02", 1189 => X"52",
        1190 => X"02", 1191 => X"53",
        1192 => X"02", 1193 => X"54",
        1194 => X"02", 1195 => X"55",
        1196 => X"02", 1197 => X"56",
        1198 => X"02", 1199 => X"57",
        1200 => X"02", 1201 => X"58",
        1202 => X"02", 1203 => X"59",
        1204 => X"02", 1205 => X"5A",
        1206 => X"02", 1207 => X"5B",
        1208 => X"02", 1209 => X"5C",
        1210 => X"02", 1211 => X"5D",
        1212 => X"02", 1213 => X"5E",
        1214 => X"02", 1215 => X"5F",
        1216 => X"02", 1217 => X"60",
        1218 => X"02", 1219 => X"61",
        1220 => X"02", 1221 => X"62",
        1222 => X"02", 1223 => X"63",
        1224 => X"02", 1225 => X"64",
        1226 => X"02", 1227 => X"65",
        1228 => X"02", 1229 => X"66",
        1230 => X"02", 1231 => X"67",
        1232 => X"02", 1233 => X"68",
        1234 => X"02", 1235 => X"69",
        1236 => X"02", 1237 => X"6A",
        1238 => X"02", 1239 => X"6B",
        1240 => X"02", 1241 => X"6C",
        1242 => X"02", 1243 => X"6D",
        1244 => X"02", 1245 => X"6E",
        1246 => X"02", 1247 => X"6F",
        1248 => X"02", 1249 => X"70",
        1250 => X"02", 1251 => X"71",
        1252 => X"02", 1253 => X"72",
        1254 => X"02", 1255 => X"73",
        1256 => X"02", 1257 => X"74",
        1258 => X"02", 1259 => X"75",
        1260 => X"02", 1261 => X"76",
        1262 => X"02", 1263 => X"77",
        1264 => X"02", 1265 => X"78",
        1266 => X"02", 1267 => X"79",
        1268 => X"02", 1269 => X"7A",
        1270 => X"02", 1271 => X"7B",
        1272 => X"02", 1273 => X"7C",
        1274 => X"02", 1275 => X"7D",
        1276 => X"02", 1277 => X"7E",
        1278 => X"02", 1279 => X"7F",
        1280 => X"02", 1281 => X"80",
        1282 => X"02", 1283 => X"81",
        1284 => X"02", 1285 => X"82",
        1286 => X"02", 1287 => X"83",
        1288 => X"02", 1289 => X"84",
        1290 => X"02", 1291 => X"85",
        1292 => X"02", 1293 => X"86",
        1294 => X"02", 1295 => X"87",
        1296 => X"02", 1297 => X"88",
        1298 => X"02", 1299 => X"89",
        1300 => X"02", 1301 => X"8A",
        1302 => X"02", 1303 => X"8B",
        1304 => X"02", 1305 => X"8C",
        1306 => X"02", 1307 => X"8D",
        1308 => X"02", 1309 => X"8E",
        1310 => X"02", 1311 => X"8F",
        1312 => X"02", 1313 => X"90",
        1314 => X"02", 1315 => X"91",
        1316 => X"02", 1317 => X"92",
        1318 => X"02", 1319 => X"93",
        1320 => X"02", 1321 => X"94",
        1322 => X"02", 1323 => X"95",
        1324 => X"02", 1325 => X"96",
        1326 => X"02", 1327 => X"97",
        1328 => X"02", 1329 => X"98",
        1330 => X"02", 1331 => X"99",
        1332 => X"02", 1333 => X"9A",
        1334 => X"02", 1335 => X"9B",
        1336 => X"02", 1337 => X"9C",
        1338 => X"02", 1339 => X"9D",
        1340 => X"02", 1341 => X"9E",
        1342 => X"02", 1343 => X"9F",
        1344 => X"02", 1345 => X"A0",
        1346 => X"02", 1347 => X"A1",
        1348 => X"02", 1349 => X"A2",
        1350 => X"02", 1351 => X"A3",
        1352 => X"02", 1353 => X"A4",
        1354 => X"02", 1355 => X"A5",
        1356 => X"02", 1357 => X"A6",
        1358 => X"02", 1359 => X"A7",
        1360 => X"02", 1361 => X"A8",
        1362 => X"02", 1363 => X"A9",
        1364 => X"02", 1365 => X"AA",
        1366 => X"02", 1367 => X"AB",
        1368 => X"02", 1369 => X"AC",
        1370 => X"02", 1371 => X"AD",
        1372 => X"02", 1373 => X"AE",
        1374 => X"02", 1375 => X"AF",
        1376 => X"02", 1377 => X"B0",
        1378 => X"02", 1379 => X"B1",
        1380 => X"02", 1381 => X"B2",
        1382 => X"02", 1383 => X"B3",
        1384 => X"02", 1385 => X"B4",
        1386 => X"02", 1387 => X"B5",
        1388 => X"02", 1389 => X"B6",
        1390 => X"02", 1391 => X"B7",
        1392 => X"02", 1393 => X"B8",
        1394 => X"02", 1395 => X"B9",
        1396 => X"02", 1397 => X"BA",
        1398 => X"02", 1399 => X"BB",
        1400 => X"02", 1401 => X"BC",
        1402 => X"02", 1403 => X"BD",
        1404 => X"02", 1405 => X"BE",
        1406 => X"02", 1407 => X"BF",
        1408 => X"02", 1409 => X"C0",
        1410 => X"02", 1411 => X"C1",
        1412 => X"02", 1413 => X"C2",
        1414 => X"02", 1415 => X"C3",
        1416 => X"02", 1417 => X"C4",
        1418 => X"02", 1419 => X"C5",
        1420 => X"02", 1421 => X"C6",
        1422 => X"02", 1423 => X"C7",
        1424 => X"02", 1425 => X"C8",
        1426 => X"02", 1427 => X"C9",
        1428 => X"02", 1429 => X"CA",
        1430 => X"02", 1431 => X"CB",
        1432 => X"02", 1433 => X"CC",
        1434 => X"02", 1435 => X"CD",
        1436 => X"02", 1437 => X"CE",
        1438 => X"02", 1439 => X"CF",
        1440 => X"02", 1441 => X"D0",
        1442 => X"02", 1443 => X"D1",
        1444 => X"02", 1445 => X"D2",
        1446 => X"02", 1447 => X"D3",
        1448 => X"02", 1449 => X"D4",
        1450 => X"02", 1451 => X"D5",
        1452 => X"02", 1453 => X"D6",
        1454 => X"02", 1455 => X"D7",
        1456 => X"02", 1457 => X"D8",
        1458 => X"02", 1459 => X"D9",
        1460 => X"02", 1461 => X"DA",
        1462 => X"02", 1463 => X"DB",
        1464 => X"02", 1465 => X"DC",
        1466 => X"02", 1467 => X"DD",
        1468 => X"02", 1469 => X"DE",
        1470 => X"02", 1471 => X"DF",
        1472 => X"02", 1473 => X"E0",
        1474 => X"02", 1475 => X"E1",
        1476 => X"02", 1477 => X"E2",
        1478 => X"02", 1479 => X"E3",
        1480 => X"02", 1481 => X"E4",
        1482 => X"02", 1483 => X"E5",
        1484 => X"02", 1485 => X"E6",
        1486 => X"02", 1487 => X"E7",
        1488 => X"02", 1489 => X"E8",
        1490 => X"02", 1491 => X"E9",
        1492 => X"02", 1493 => X"EA",
        1494 => X"02", 1495 => X"EB",
        1496 => X"02", 1497 => X"EC",
        1498 => X"02", 1499 => X"ED"
    )
);
    
BEGIN

    project_cmp : project_io PORT MAP (
        clk => clk,
        rst => rst,
        enable => enable,
        done => done,
        in_read_enable => in_read_enable,
        in_index => in_index,
        in_data => in_data,
        out_write_enable => out_write_enable,
        out_index => out_index,
        out_data => out_data,
        in_buff_size => in_buff_size,
        out_buff_size => out_buff_size
    );

    p_clock : PROCESS 
    BEGIN 
        clk <= '0';
        wait for 10 ns;
        clk <= '1';
        wait for 10 ns;
    END PROCESS p_clock;


    process
    begin
        wait for 60100 ns;
        report "end" severity failure;
    end process;

    PROCESS (clk)
    begin
        if rising_edge(clk) then
            if done = '1' then
                enable <= not done;
                
            elsif enable = '0' then
                if curr_buffer = BUFFER_NUM then
                    report "end" severity failure;
                end if;
                in_ram <= buffer_array(curr_buffer);

                curr_buffer <= curr_buffer + 1;

                enable <= '1';
            end if;
        end if;

    end process;
    

    p_ram_reader : PROCESS (clk)
BEGIN 
    IF rising_edge(clk) AND enable = '1' AND in_read_enable = '1' THEN
        IF in_index >= 0 AND in_index <= IN_RAM_SIZE - 1 THEN
            in_data <= in_ram(in_index);
        ELSE
            report "Invalid in_index: " & integer'image(in_index) severity warning;
            in_data <= (others => '0'); -- assign a safe default
        END IF;
    END IF;
END PROCESS p_ram_reader;


    p_ram_output : PROCESS (clk)
    variable line_out : line;
    BEGIN 
        IF rising_edge(clk) AND out_write_enable = '1' AND enable = '1' THEN
            
            write (line_out, to_integer(unsigned(out_data)));
            writeline (output, line_out);
        END IF;
    END PROCESS p_ram_output;

    

END architecture behavioural;
